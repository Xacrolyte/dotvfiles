version https://git-lfs.github.com/spec/v1
oid sha256:c6e95305eb526ec7f40c8018783f5adf9a36d03c2b91b3a2313a8c2da17ab9b9
size 2984
